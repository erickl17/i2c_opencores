package i2c_env_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import wishbone_agent_pkg::*;

  `include "i2c_env_cfg.svh"
  `include "i2c_env.svh"
endpackage : i2c_env_pkg